library verilog;
use verilog.vl_types.all;
entity DECODE2_4_vlg_vec_tst is
end DECODE2_4_vlg_vec_tst;
