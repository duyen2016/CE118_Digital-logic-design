library verilog;
use verilog.vl_types.all;
entity PRCS_vlg_vec_tst is
end PRCS_vlg_vec_tst;
