library verilog;
use verilog.vl_types.all;
entity DECODE2_4_vlg_check_tst is
    port(
        D               : in     vl_logic_vector(3 downto 0);
        sampler_rx      : in     vl_logic
    );
end DECODE2_4_vlg_check_tst;
