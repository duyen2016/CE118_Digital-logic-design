library verilog;
use verilog.vl_types.all;
entity MEALY_LBSMSSV_vlg_vec_tst is
end MEALY_LBSMSSV_vlg_vec_tst;
