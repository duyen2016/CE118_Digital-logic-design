library verilog;
use verilog.vl_types.all;
entity MEALY_LBSMSSV_vlg_check_tst is
    port(
        OUTPUT          : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end MEALY_LBSMSSV_vlg_check_tst;
