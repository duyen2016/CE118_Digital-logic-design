library verilog;
use verilog.vl_types.all;
entity RAM4x8bit_vlg_vec_tst is
end RAM4x8bit_vlg_vec_tst;
