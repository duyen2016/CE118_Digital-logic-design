library verilog;
use verilog.vl_types.all;
entity PRSC_DE2KIT_vlg_vec_tst is
end PRSC_DE2KIT_vlg_vec_tst;
