library verilog;
use verilog.vl_types.all;
entity RAM16x8bit_vlg_vec_tst is
end RAM16x8bit_vlg_vec_tst;
