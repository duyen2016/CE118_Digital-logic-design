library verilog;
use verilog.vl_types.all;
entity MEALY_MSSV_vlg_vec_tst is
end MEALY_MSSV_vlg_vec_tst;
