library verilog;
use verilog.vl_types.all;
entity MOORE_MSSV_vlg_vec_tst is
end MOORE_MSSV_vlg_vec_tst;
