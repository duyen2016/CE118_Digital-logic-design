library verilog;
use verilog.vl_types.all;
entity RAM32x8bit_vlg_vec_tst is
end RAM32x8bit_vlg_vec_tst;
