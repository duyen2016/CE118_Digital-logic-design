library verilog;
use verilog.vl_types.all;
entity CONTROL_vlg_vec_tst is
end CONTROL_vlg_vec_tst;
