library verilog;
use verilog.vl_types.all;
entity MC_vlg_vec_tst is
end MC_vlg_vec_tst;
