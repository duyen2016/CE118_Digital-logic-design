library verilog;
use verilog.vl_types.all;
entity NHAN4BIT_vlg_vec_tst is
end NHAN4BIT_vlg_vec_tst;
