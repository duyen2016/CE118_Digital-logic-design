library verilog;
use verilog.vl_types.all;
entity LU_vlg_vec_tst is
end LU_vlg_vec_tst;
